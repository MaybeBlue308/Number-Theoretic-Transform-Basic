
module rom_zeta(
 //   input wire clk,
    input  wire [6:0]  addr,
    output reg  [11:0] data
);
    reg [11:0] rom [0:127];
    initial begin
 rom[0]  = 12'h001;
        rom[1]  = 12'h6C1;
        rom[2]  = 12'hA14;
        rom[3]  = 12'hCD9;
        rom[4]  = 12'hA52;
        rom[5]  = 12'h276;
        rom[6]  = 12'h769;
        rom[7]  = 12'h350;
        rom[8]  = 12'h426;
        rom[9]  = 12'h77F;
        rom[10] = 12'h0C1;
        rom[11] = 12'h31D;
        rom[12] = 12'hAE2;
        rom[13] = 12'hCBC;
        rom[14] = 12'h239;
        rom[15] = 12'h6D2;
        rom[16] = 12'h128;
        rom[17] = 12'h98F;
        rom[18] = 12'h53B;
        rom[19] = 12'h5C4;
        rom[20] = 12'hBE6;
        rom[21] = 12'h038;
        rom[22] = 12'h8C0;
        rom[23] = 12'h535;
        rom[24] = 12'h592;
        rom[25] = 12'h82E;
        rom[26] = 12'h217;
        rom[27] = 12'hB42;
        rom[28] = 12'h959;
        rom[29] = 12'hB3F;
        rom[30] = 12'h7B6;
        rom[31] = 12'h335;
        rom[32] = 12'h121;
        rom[33] = 12'h14B;
        rom[34] = 12'hCB5;
        rom[35] = 12'h6DC;
        rom[36] = 12'h4AD;
        rom[37] = 12'h900;
        rom[38] = 12'h8E5;
        rom[39] = 12'h807;
        rom[40] = 12'h28A;
        rom[41] = 12'h7B9;
        rom[42] = 12'h9D1;
        rom[43] = 12'h278;
        rom[44] = 12'hB31;
        rom[45] = 12'h021;
        rom[46] = 12'h528;
        rom[47] = 12'h77B;
        rom[48] = 12'h90F;
        rom[49] = 12'h59B;
        rom[50] = 12'h327;
        rom[51] = 12'h1C4;
        rom[52] = 12'h59E;
        rom[53] = 12'hB34;
        rom[54] = 12'h5FE;
        rom[55] = 12'h962;
        rom[56] = 12'hA57;
        rom[57] = 12'hA39;
        rom[58] = 12'h5C9;
        rom[59] = 12'h288;
        rom[60] = 12'h9AA;
        rom[61] = 12'hC26;
        rom[62] = 12'h4CB;
        rom[63] = 12'h38E;
        rom[64] = 12'h011;
        rom[65] = 12'hAC9;
        rom[66] = 12'h247;
        rom[67] = 12'hA59;
        rom[68] = 12'h665;
        rom[69] = 12'h2D3;
        rom[70] = 12'h8F0;
        rom[71] = 12'h44C;
        rom[72] = 12'h581;
        rom[73] = 12'hA66;
        rom[74] = 12'hCD1;
        rom[75] = 12'h0E9;
        rom[76] = 12'h2F4;
        rom[77] = 12'h86C;
        rom[78] = 12'hBC7;
        rom[79] = 12'hBEA;
        rom[80] = 12'h6A7;
        rom[81] = 12'h673;
        rom[82] = 12'hAE5;
        rom[83] = 12'h6FD;
        rom[84] = 12'h737;
        rom[85] = 12'h3B8;
        rom[86] = 12'h5B5;
        rom[87] = 12'hA7F;
        rom[88] = 12'h3AB;
        rom[89] = 12'h904;
        rom[90] = 12'h985;
        rom[91] = 12'h954;
        rom[92] = 12'h2DD;
        rom[93] = 12'h921;
        rom[94] = 12'h10C;
        rom[95] = 12'h281;
        rom[96] = 12'h630;
        rom[97] = 12'h8FA;
        rom[98] = 12'h7F5;
        rom[99] = 12'hC94;
        rom[100]= 12'h177;
        rom[101]= 12'h9F5;
        rom[102]= 12'h82A;
        rom[103]= 12'h66D;
        rom[104]= 12'h427;
        rom[105]= 12'h13F;
        rom[106]= 12'hAD5;
        rom[107]= 12'h2F5;
        rom[108]= 12'h833;
        rom[109]= 12'h231;
        rom[110]= 12'h9A2;
        rom[111]= 12'hA22;
        rom[112]= 12'hAF4;
        rom[113]= 12'h444;
        rom[114]= 12'h193;
        rom[115]= 12'h402;
        rom[116]= 12'h477;
        rom[117]= 12'h866;
        rom[118]= 12'hAD7;
        rom[119]= 12'h376;
        rom[120]= 12'h6BA;
        rom[121]= 12'h4BC;
        rom[122]= 12'h752;
        rom[123]= 12'h405;
        rom[124]= 12'h83E;
        rom[125]= 12'hB77;
        rom[126]= 12'h375;
        rom[127]= 12'h86A;
    end
    always @(*) begin
        data = rom[addr];
    end
endmodule


